module add16(
    input [7:0] a, b,
    output [15:0] sum
);
endmodule